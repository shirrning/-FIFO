`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/07/22 20:28:21
// Design Name: 
// Module Name: yasuo3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module     yasuo3(j000,j100,j200,j20_s,j20_c);

input   [23:0] j000,j100;
input   [22:0] j200;

output  [28:0] j20_s;
output  [26:0] j20_c;

wire    [28:0] j20_s;
wire    [26:0] j20_c;


assign j20_s[28]=j200[19];
assign j20_s[3]=j000[3];
assign j20_s[2]=j000[2];
assign j20_s[1]=j000[1];
assign j20_s[0]=j000[0];
assign j20_c[26]=j200[22];
assign j20_c[25]=j200[21];
assign j20_c[24]=j200[20];

add3  a1 (.a(1'b0),     .b(j100[23]), .c(j200[18]), .si(j20_s[27]), .ci(j20_c[23]));
add3  a2 (.a(1'b0),     .b(j100[22]), .c(j200[17]), .si(j20_s[26]), .ci(j20_c[22]));
add3  a3 (.a(1'b0),     .b(j100[21]), .c(j200[16]), .si(j20_s[25]), .ci(j20_c[21]));
add3  a4 (.a(1'b0),     .b(j100[20]), .c(j200[15]), .si(j20_s[24]), .ci(j20_c[20]));
add3  a5 (.a(j000[23]), .b(j100[19]), .c(j200[14]), .si(j20_s[23]), .ci(j20_c[19]));
add3  a6 (.a(j000[22]), .b(j100[18]), .c(j200[13]), .si(j20_s[22]), .ci(j20_c[18]));
add3  a7 (.a(j000[21]), .b(j100[17]), .c(j200[12]), .si(j20_s[21]), .ci(j20_c[17]));
add3  a8 (.a(j000[20]), .b(j100[16]), .c(j200[11]), .si(j20_s[20]), .ci(j20_c[16]));
add3  a9 (.a(j000[19]), .b(j100[15]), .c(j200[10]), .si(j20_s[19]), .ci(j20_c[15]));
add3  a10(.a(j000[18]), .b(j100[14]), .c(j200[9]),  .si(j20_s[18]), .ci(j20_c[14]));
add3  a11(.a(j000[17]), .b(j100[13]), .c(j200[8]),  .si(j20_s[17]), .ci(j20_c[13]));
add3  a12(.a(j000[16]), .b(j100[12]), .c(j200[7]),  .si(j20_s[16]), .ci(j20_c[12]));
add3  a13(.a(j000[15]), .b(j100[11]), .c(j200[6]),  .si(j20_s[15]), .ci(j20_c[11]));
add3  a14(.a(j000[14]), .b(j100[10]), .c(j200[5]),  .si(j20_s[14]), .ci(j20_c[10]));
add3  a15(.a(j000[13]), .b(j100[9]),  .c(j200[4]),  .si(j20_s[13]), .ci(j20_c[9]));
add3  a16(.a(j000[12]), .b(j100[8]),  .c(j200[3]),  .si(j20_s[12]), .ci(j20_c[8]));
add3  a17(.a(j000[11]), .b(j100[7]),  .c(j200[2]),  .si(j20_s[11]), .ci(j20_c[7]));
add3  a18(.a(j000[10]), .b(j100[6]),  .c(j200[1]),  .si(j20_s[10]), .ci(j20_c[6]));
add3  a19(.a(j000[9]),  .b(j100[5]),  .c(j200[0]),  .si(j20_s[9]),  .ci(j20_c[5]));
add3  a20(.a(j000[8]),  .b(j100[4]),  .c(1'b0),     .si(j20_s[8]),  .ci(j20_c[4]));
add3  a21(.a(j000[7]),  .b(j100[3]),  .c(1'b0),     .si(j20_s[7]),  .ci(j20_c[3]));
add3  a22(.a(j000[6]),  .b(j100[2]),  .c(1'b0),     .si(j20_s[6]),  .ci(j20_c[2]));
add3  a23(.a(j000[5]),  .b(j100[1]),  .c(1'b0),     .si(j20_s[5]),  .ci(j20_c[1]));
add3  a24(.a(j000[4]),  .b(j100[0]),  .c(1'b0),     .si(j20_s[4]),  .ci(j20_c[0]));

endmodule

