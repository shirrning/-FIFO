`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/07/22 20:28:21
// Design Name: 
// Module Name: yasuo1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module     yasuo1(j0,j1,j2,j3,j4,j5,j6,j7,j8,j0_s,j0_c,j1_s,j1_c,j2_s,j2_c);

input    [19:0] j0;
input    [18:0] j1,j2,j3,j4,j5,j6;
input    [17:0] j7;
input    [16:0] j8; 

output   [21:0] j0_s,j1_s;
output   [19:0] j0_c,j1_c,j2_s;
output   [17:0] j2_c;

wire     [21:0] j0_s,j1_s;
wire     [19:0] j0_c,j1_c,j2_s;
wire     [17:0] j2_c;

//j0_s,j0_c

assign j0_s[21]=j2[17];
assign j0_s[1]=j0[1];
assign j0_s[0]=j0[0];
assign j0_c[19]=j2[18];

add3  a1 (.a(1'b0), .b(j1[18]), .c(j2[16]), .si(j0_s[20]), .ci(j0_c[18]));
add3  a2 (.a(j0[19]), .b(j1[17]), .c(j2[15]), .si(j0_s[19]), .ci(j0_c[17]));
add3  a3 (.a(j0[18]), .b(j1[16]), .c(j2[14]), .si(j0_s[18]), .ci(j0_c[16]));
add3  a4 (.a(j0[17]), .b(j1[15]), .c(j2[13]), .si(j0_s[17]), .ci(j0_c[15]));
add3  a5 (.a(j0[16]), .b(j1[14]), .c(j2[12]), .si(j0_s[16]), .ci(j0_c[14]));
add3  a6 (.a(j0[15]), .b(j1[13]), .c(j2[11]), .si(j0_s[15]), .ci(j0_c[13]));
add3  a7 (.a(j0[14]), .b(j1[12]), .c(j2[10]), .si(j0_s[14]), .ci(j0_c[12]));
add3  a8 (.a(j0[13]), .b(j1[11]), .c(j2[9]),  .si(j0_s[13]), .ci(j0_c[11]));
add3  a9 (.a(j0[12]), .b(j1[10]), .c(j2[8]),  .si(j0_s[12]), .ci(j0_c[10]));
add3  a10(.a(j0[11]), .b(j1[9]),  .c(j2[7]),  .si(j0_s[11]), .ci(j0_c[9]));
add3  a11(.a(j0[10]), .b(j1[8]),  .c(j2[6]),  .si(j0_s[10]), .ci(j0_c[8]));
add3  a12(.a(j0[9]),  .b(j1[7]),  .c(j2[5]),  .si(j0_s[9]),  .ci(j0_c[7]));
add3  a13(.a(j0[8]),  .b(j1[6]),  .c(j2[4]),  .si(j0_s[8]),  .ci(j0_c[6]));
add3  a14(.a(j0[7]),  .b(j1[5]),  .c(j2[3]),  .si(j0_s[7]),  .ci(j0_c[5]));
add3  a15(.a(j0[6]),  .b(j1[4]),  .c(j2[2]),  .si(j0_s[6]),  .ci(j0_c[4]));
add3  a16(.a(j0[5]),  .b(j1[3]),  .c(j2[1]),  .si(j0_s[5]),  .ci(j0_c[3]));
add3  a17(.a(j0[4]),  .b(j1[2]),  .c(j2[0]),  .si(j0_s[4]),  .ci(j0_c[2]));
add3  a18(.a(j0[3]),  .b(j1[1]),  .c(1'b0),     .si(j0_s[3]),  .ci(j0_c[1]));
add3  a19(.a(j0[2]),  .b(j1[0]),  .c(1'b0),     .si(j0_s[2]),  .ci(j0_c[0]));



//j1_s,j1_c


assign j1_s[21]=j5[17];
assign j1_s[1]=j3[1];
assign j1_s[0]=j3[0];
assign j1_c[19]=j5[18];

add3  a20(.a(1'b0), .b(j4[18]), .c(j5[16]), .si(j1_s[20]), .ci(j1_c[18]));
add3  a21(.a(1'b0), .b(j4[17]), .c(j5[15]), .si(j1_s[19]), .ci(j1_c[17]));
add3  a22(.a(j3[18]), .b(j4[16]), .c(j5[14]), .si(j1_s[18]), .ci(j1_c[16]));
add3  a23(.a(j3[17]), .b(j4[15]), .c(j5[13]), .si(j1_s[17]), .ci(j1_c[15]));
add3  a24(.a(j3[16]), .b(j4[14]), .c(j5[12]), .si(j1_s[16]), .ci(j1_c[14]));
add3  a25(.a(j3[15]), .b(j4[13]), .c(j5[11]), .si(j1_s[15]), .ci(j1_c[13]));
add3  a26(.a(j3[14]), .b(j4[12]), .c(j5[10]), .si(j1_s[14]), .ci(j1_c[12]));
add3  a27(.a(j3[13]), .b(j4[11]), .c(j5[9]),  .si(j1_s[13]), .ci(j1_c[11]));
add3  a28(.a(j3[12]), .b(j4[10]), .c(j5[8]),  .si(j1_s[12]), .ci(j1_c[10]));
add3  a29(.a(j3[11]), .b(j4[9]),  .c(j5[7]),  .si(j1_s[11]), .ci(j1_c[9]));
add3  a30(.a(j3[10]), .b(j4[8]),  .c(j5[6]),  .si(j1_s[10]), .ci(j1_c[8]));
add3  a31(.a(j3[9]),  .b(j4[7]),  .c(j5[5]),  .si(j1_s[9]),  .ci(j1_c[7]));
add3  a32(.a(j3[8]),  .b(j4[6]),  .c(j5[4]),  .si(j1_s[8]),  .ci(j1_c[6]));
add3  a33(.a(j3[7]),  .b(j4[5]),  .c(j5[3]),  .si(j1_s[7]),  .ci(j1_c[5]));
add3  a34(.a(j3[6]),  .b(j4[4]),  .c(j5[2]),  .si(j1_s[6]),  .ci(j1_c[4]));
add3  a35(.a(j3[5]),  .b(j4[3]),  .c(j5[1]),  .si(j1_s[5]),  .ci(j1_c[3]));
add3  a36(.a(j3[4]),  .b(j4[2]),  .c(j5[0]),  .si(j1_s[4]),  .ci(j1_c[2]));
add3  a37(.a(j3[3]),  .b(j4[1]),  .c(1'b0),     .si(j1_s[3]),  .ci(j1_c[1]));
add3  a38(.a(j3[2]),  .b(j4[0]),  .c(1'b0),     .si(j1_s[2]),  .ci(j1_c[0]));

//j2_s,j2_c

assign j2_s[1]=j6[1];
assign j2_s[0]=j6[0];

add3  a39(.a(1'b0), .b(j7[17]), .c(j8[15]), .si(j2_s[19]), .ci(j2_c[17]));
add3  a40(.a(j6[18]), .b(j7[16]), .c(j8[14]), .si(j2_s[18]), .ci(j2_c[16]));
add3  a41(.a(j6[17]), .b(j7[15]), .c(j8[13]), .si(j2_s[17]), .ci(j2_c[15]));
add3  a42(.a(j6[16]), .b(j7[14]), .c(j8[12]), .si(j2_s[16]), .ci(j2_c[14]));
add3  a43(.a(j6[15]), .b(j7[13]), .c(j8[11]), .si(j2_s[15]), .ci(j2_c[13]));
add3  a44(.a(j6[14]), .b(j7[12]), .c(j8[10]), .si(j2_s[14]), .ci(j2_c[12]));
add3  a45(.a(j6[13]), .b(j7[11]), .c(j8[9]),  .si(j2_s[13]), .ci(j2_c[11]));
add3  a46(.a(j6[12]), .b(j7[10]), .c(j8[8]),  .si(j2_s[12]), .ci(j2_c[10]));
add3  a47(.a(j6[11]), .b(j7[9]),  .c(j8[7]),  .si(j2_s[11]), .ci(j2_c[9]));
add3  a48(.a(j6[10]), .b(j7[8]),  .c(j8[6]),  .si(j2_s[10]), .ci(j2_c[8]));
add3  a49(.a(j6[9]),  .b(j7[7]),  .c(j8[5]),  .si(j2_s[9]),  .ci(j2_c[7]));
add3  a50(.a(j6[8]),  .b(j7[6]),  .c(j8[4]),  .si(j2_s[8]),  .ci(j2_c[6]));
add3  a51(.a(j6[7]),  .b(j7[5]),  .c(j8[3]),  .si(j2_s[7]),  .ci(j2_c[5]));
add3  a52(.a(j6[6]),  .b(j7[4]),  .c(j8[2]),  .si(j2_s[6]),  .ci(j2_c[4]));
add3  a53(.a(j6[5]),  .b(j7[3]),  .c(j8[1]),  .si(j2_s[5]),  .ci(j2_c[3]));
add3  a54(.a(j6[4]),  .b(j7[2]),  .c(j8[0]),  .si(j2_s[4]),  .ci(j2_c[2]));
add3  a55(.a(j6[3]),  .b(j7[1]),  .c(1'b0),     .si(j2_s[3]),  .ci(j2_c[1]));
add3  a56(.a(j6[2]),  .b(j7[0]),  .c(1'b0),     .si(j2_s[2]),  .ci(j2_c[0]));

endmodule
