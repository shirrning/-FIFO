`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/07/22 20:28:21
// Design Name: 
// Module Name: yasuo4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module     yasuo4(j10,j20,j30,j0000,j1000);

input   [28:0] j10;
input   [26:0] j20;
input   [19:0] j30;
output  [31:0] j0000;
output  [26:0] j1000;

wire    [31:0] j0000;
wire    [26:0] j1000;

assign j0000[4]=j10[4];
assign j0000[3]=j10[3];
assign j0000[2]=j10[2];
assign j0000[1]=j10[1];
assign j0000[0]=j10[0];


add3  a1 (.a(1'b0),    .b(j20[26]), .c(j30[18]), .si(j0000[31]), .ci(j1000[26]));
add3  a2 (.a(1'b0),    .b(j20[25]), .c(j30[17]), .si(j0000[30]), .ci(j1000[25]));
add3  a3 (.a(1'b0),    .b(j20[24]), .c(j30[16]), .si(j0000[29]), .ci(j1000[24]));
add3  a4 (.a(j10[28]), .b(j20[23]), .c(j30[15]), .si(j0000[28]), .ci(j1000[23]));
add3  a5 (.a(j10[27]), .b(j20[22]), .c(j30[14]), .si(j0000[27]), .ci(j1000[22]));
add3  a6 (.a(j10[26]), .b(j20[21]), .c(j30[13]), .si(j0000[26]), .ci(j1000[21]));
add3  a7 (.a(j10[25]), .b(j20[20]), .c(j30[12]), .si(j0000[25]), .ci(j1000[20]));
add3  a8 (.a(j10[24]), .b(j20[19]), .c(j30[11]), .si(j0000[24]), .ci(j1000[19]));
add3  a9 (.a(j10[23]), .b(j20[18]), .c(j30[10]), .si(j0000[23]), .ci(j1000[18]));
add3  a10(.a(j10[22]), .b(j20[17]), .c(j30[9]),  .si(j0000[22]), .ci(j1000[17]));
add3  a11(.a(j10[21]), .b(j20[16]), .c(j30[8]),  .si(j0000[21]), .ci(j1000[16]));
add3  a12(.a(j10[20]), .b(j20[15]), .c(j30[7]),  .si(j0000[20]), .ci(j1000[15]));
add3  a13(.a(j10[19]), .b(j20[14]), .c(j30[6]),  .si(j0000[19]), .ci(j1000[14]));
add3  a14(.a(j10[18]), .b(j20[13]), .c(j30[5]),  .si(j0000[18]), .ci(j1000[13]));
add3  a15(.a(j10[17]), .b(j20[12]), .c(j30[4]),  .si(j0000[17]), .ci(j1000[12]));
add3  a16(.a(j10[16]), .b(j20[11]), .c(j30[3]),  .si(j0000[16]), .ci(j1000[11]));
add3  a17(.a(j10[15]), .b(j20[10]), .c(j30[2]),  .si(j0000[15]), .ci(j1000[10]));
add3  a18(.a(j10[14]), .b(j20[9]),  .c(j30[1]),  .si(j0000[14]), .ci(j1000[9]));
add3  a19(.a(j10[13]), .b(j20[8]),  .c(j30[0]),  .si(j0000[13]), .ci(j1000[8]));
add3  a20(.a(j10[12]), .b(j20[7]),  .c(1'b0),    .si(j0000[12]), .ci(j1000[7]));
add3  a21(.a(j10[11]), .b(j20[6]),  .c(1'b0),    .si(j0000[11]), .ci(j1000[6]));
add3  a22(.a(j10[10]), .b(j20[5]),  .c(1'b0),    .si(j0000[10]), .ci(j1000[5]));
add3  a23(.a(j10[9]),  .b(j20[4]),  .c(1'b0),    .si(j0000[9]),  .ci(j1000[4]));
add3  a24(.a(j10[8]),  .b(j20[3]),  .c(1'b0),    .si(j0000[8]),  .ci(j1000[3]));
add3  a25(.a(j10[7]),  .b(j20[2]),  .c(1'b0),    .si(j0000[7]),  .ci(j1000[2]));
add3  a26(.a(j10[6]),  .b(j20[1]),  .c(1'b0),    .si(j0000[6]),  .ci(j1000[1]));
add3  a27(.a(j10[5]),  .b(j20[0]),  .c(1'b0),    .si(j0000[5]),  .ci(j1000[0]));

endmodule
